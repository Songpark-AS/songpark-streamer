----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 06/15/2019 04:04:36 PM
-- Design Name: 
-- Module Name: RTLTD_SLV_PIPELINE_SEARCH - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity RTLTD_SLV_PIPELINE_SEARCH is
--  Port ( );
end RTLTD_SLV_PIPELINE_SEARCH;

architecture Behavioral of RTLTD_SLV_PIPELINE_SEARCH is

begin


end Behavioral;
