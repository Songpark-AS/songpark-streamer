----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 08/27/2020 08:46:06 PM
-- Design Name: 
-- Module Name: pck_interpolator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package pck_interpolator is

    attribute enum_encoding: string;

--    function stdl (arg: boolean) return std_logic;

--    function stdl (arg: integer) return std_logic;

--    function to_unsigned (arg: boolean; size: natural) return unsigned;

--    function to_signed (arg: boolean; size: natural) return signed;

--    function to_integer(arg: boolean) return integer;

--    function to_integer(arg: std_logic) return integer;

--    function to_unsigned (arg: std_logic; size: natural) return unsigned;

--    function to_signed (arg: std_logic; size: natural) return signed;

    function bool (arg: std_logic) return boolean;

    function bool (arg: unsigned) return boolean;

    function bool (arg: signed) return boolean;

    function bool (arg: integer) return boolean;

    function "-" (arg: unsigned) return signed;

    function tern_op(cond: boolean; if_true: std_logic; if_false: std_logic) return std_logic;

    function tern_op(cond: boolean; if_true: unsigned; if_false: unsigned) return unsigned;

    function tern_op(cond: boolean; if_true: signed; if_false: signed) return signed;

end pck_interpolator;


package body pck_interpolator is

    function stdl (arg: boolean) return std_logic is
    begin
        if arg then
            return '1';
        else
            return '0';
        end if;
    end function stdl;

    function stdl (arg: integer) return std_logic is
    begin
        if arg /= 0 then
            return '1';
        else
            return '0';
        end if;
    end function stdl;


--    function to_unsigned (arg: boolean; size: natural) return unsigned is
--        variable res: unsigned(size-1 downto 0) := (others => '0');
--    begin
--        if arg then
--            res(0):= '1';
--        end if;
--        return res;
--    end function to_unsigned;

--    function to_signed (arg: boolean; size: natural) return signed is
--        variable res: signed(size-1 downto 0) := (others => '0');
--    begin
--        if arg then
--            res(0) := '1';
--        end if;
--        return res; 
--    end function to_signed;

--    function to_integer(arg: boolean) return integer is
--    begin
--        if arg then
--            return 1;
--        else
--            return 0;
--        end if;
--    end function to_integer;

--    function to_integer(arg: std_logic) return integer is
--    begin
--        if arg = '1' then
--            return 1;
--        else
--            return 0;
--        end if;
--    end function to_integer;

--    function to_unsigned (arg: std_logic; size: natural) return unsigned is
--        variable res: unsigned(size-1 downto 0) := (others => '0');
--    begin
--        res(0):= arg;
--        return res;
--    end function to_unsigned;

--    function to_signed (arg: std_logic; size: natural) return signed is
--        variable res: signed(size-1 downto 0) := (others => '0');
--    begin
--        res(0) := arg;
--        return res; 
--    end function to_signed;

    function bool (arg: std_logic) return boolean is
    begin
        return arg = '1';
    end function bool;

    function bool (arg: unsigned) return boolean is
    begin
        return arg /= 0;
    end function bool;

    function bool (arg: signed) return boolean is
    begin
        return arg /= 0;
    end function bool;

    function bool (arg: integer) return boolean is
    begin
        return arg /= 0;
    end function bool;

    function "-" (arg: unsigned) return signed is
    begin
        return - signed(resize(arg, arg'length+1));
    end function "-";

    function tern_op(cond: boolean; if_true: std_logic; if_false: std_logic) return std_logic is
    begin
        if cond then
            return if_true;
        else
            return if_false;
        end if;
    end function tern_op;

    function tern_op(cond: boolean; if_true: unsigned; if_false: unsigned) return unsigned is
    begin
        if cond then
            return if_true;
        else
            return if_false;
        end if;
    end function tern_op;

    function tern_op(cond: boolean; if_true: signed; if_false: signed) return signed is
    begin
        if cond then
            return if_true;
        else
            return if_false;
        end if;
    end function tern_op;

end pck_interpolator;